module Simple_counter_switch_fpga(
								input clk,
								output reg [0:7]d	
												);

endmodule 

